
`timescale 1 ns / 1 ps

/**
 * @note:
 * 1. size of image must be integral multiple of C_M_AXI_DATA_WIDTH * C_M_AXI_BURST_LEN.
 * 2. the sof [start of frame] must be 1'b1 for first image data.
 * 3. width of image must be integral multiple of C_M_AXI_DATA_WIDTH.
 */
module PVDMA_M_AXI_R #
(
	// Users to add parameters here
	parameter integer C_IMG_WBITS	= 12,
	parameter integer C_IMG_HBITS	= 12,
	parameter integer C_IMG_WIDTH	= 1280,
	parameter integer C_IMG_HEIGHT	= 800,

	// User parameters ends
	// Do not modify the parameters beyond this line

	// Burst Length. Supports 1, 2, 4, 8, 16, 32, 64, 128, 256 burst lengths
	parameter integer C_M_AXI_BURST_LEN	= 16,
	// Thread ID Width
	parameter integer C_M_AXI_ID_WIDTH	= 1,
	// Width of Address Bus
	parameter integer C_M_AXI_ADDR_WIDTH	= 32,
	// Width of Data Bus
	parameter integer C_M_AXI_DATA_WIDTH	= 32
)
(
	// Users to add ports here
	output wire sof,
	output wire eol,
	output wire [C_M_AXI_DATA_WIDTH-1 : 0] dout,
	output wire wr_en,
	input wire full,

	output reg frame_pulse,
	input wire [C_M_AXI_ADDR_WIDTH-1 : 0] base_addr,

	// User ports ends
	// Do not modify the ports beyond this line

	// Global Clock Signal.
	input wire  M_AXI_ACLK,
	// Global Reset Singal. This Signal is Active Low
	input wire  M_AXI_ARESETN,

	// Master Interface Read Address.
	output wire [C_M_AXI_ID_WIDTH-1 : 0] M_AXI_ARID,
	// Read address. This signal indicates the initial
// address of a read burst transaction.
	output wire [C_M_AXI_ADDR_WIDTH-1 : 0] M_AXI_ARADDR,
	// Burst length. The burst length gives the exact number of transfers in a burst
	output wire [7 : 0] M_AXI_ARLEN,
	// Burst size. This signal indicates the size of each transfer in the burst
	output wire [2 : 0] M_AXI_ARSIZE,
	// Burst type. The burst type and the size information,
// determine how the address for each transfer within the burst is calculated.
	output wire [1 : 0] M_AXI_ARBURST,
	// Lock type. Provides additional information about the
// atomic characteristics of the transfer.
	output wire  M_AXI_ARLOCK,
	// Memory type. This signal indicates how transactions
// are required to progress through a system.
	output wire [3 : 0] M_AXI_ARCACHE,
	// Protection type. This signal indicates the privilege
// and security level of the transaction, and whether
// the transaction is a data access or an instruction access.
	output wire [2 : 0] M_AXI_ARPROT,
	// Quality of Service, QoS identifier sent for each read transaction
	output wire [3 : 0] M_AXI_ARQOS,
	// Write address valid. This signal indicates that
// the channel is signaling valid read address and control information
	output wire  M_AXI_ARVALID,
	// Read address ready. This signal indicates that
// the slave is ready to accept an address and associated control signals
	input wire  M_AXI_ARREADY,
	// Read ID tag. This signal is the identification tag
// for the read data group of signals generated by the slave.
	input wire [C_M_AXI_ID_WIDTH-1 : 0] M_AXI_RID,
	// Master Read Data
	input wire [C_M_AXI_DATA_WIDTH-1 : 0] M_AXI_RDATA,
	// Read response. This signal indicates the status of the read transfer
	input wire [1 : 0] M_AXI_RRESP,
	// Read last. This signal indicates the last transfer in a read burst
	input wire  M_AXI_RLAST,
	// Read valid. This signal indicates that the channel
// is signaling the required read data.
	input wire  M_AXI_RVALID,
	// Read ready. This signal indicates that the master can
// accept the read data and response information.
	output wire  M_AXI_RREADY
);


	// function called clogb2 that returns an integer which has the
	//value of the ceiling of the log base 2

	// function called clogb2 that returns an integer which has the
	// value of the ceiling of the log base 2.
	function integer clogb2 (input integer bit_depth);
	begin
	for(clogb2=0; bit_depth>0; clogb2=clogb2+1)
	bit_depth = bit_depth >> 1;
	end
	endfunction

	// C_TRANSACTIONS_NUM is the width of the index counter for
	// number of write or read transaction.
	localparam integer C_TRANSACTIONS_NUM = clogb2(C_M_AXI_BURST_LEN-1);

	// Burst length for transactions, in C_M_AXI_DATA_WIDTHs.
	// Non-2^n lengths will eventually cause bursts across 4K address boundaries.
	localparam integer C_MASTER_LENGTH	= 12;
	// total number of burst transfers is master length divided by burst length and burst size
	localparam integer C_NO_BURSTS_REQ = C_MASTER_LENGTH-clogb2((C_M_AXI_BURST_LEN*C_M_AXI_DATA_WIDTH/8)-1);

	// AXI4LITE signals
	//AXI4 internal temp signals
	reg [C_M_AXI_ADDR_WIDTH-1 : 0] 	axi_araddr;
	reg  	axi_arvalid;
	wire  	axi_rready;
	//read beat count in a burst
	reg [C_TRANSACTIONS_NUM : 0] 	read_index;
	//size of C_M_AXI_BURST_LEN length burst in bytes
	wire [C_TRANSACTIONS_NUM+2 : 0] 	burst_size_bytes;
	/// @note: don't across 4K edge
	reg  	start_single_burst_read;
	reg  	burst_read_active;
	//Interface response error flags
	wire  	read_resp_error;
	wire  	rnext;

	reg	r_sof;
	reg	r_eol;
	reg [C_IMG_WBITS-1 : 0] r_img_col_idx;
	reg [C_IMG_HBITS-1 : 0] r_img_row_idx;


	// I/O Connections assignments
	assign sof		= r_sof;
	assign eol		= r_eol;
	assign dout		= M_AXI_RDATA;
	assign wr_en		= rnext;
	assign axi_rready	= ~full;

	//Read Address (AR)
	assign M_AXI_ARID	= 'b0;
	assign M_AXI_ARADDR	= axi_araddr;
	//Burst LENgth is number of transaction beats, minus 1
	assign M_AXI_ARLEN	= C_M_AXI_BURST_LEN - 1;
	//Size should be C_M_AXI_DATA_WIDTH, in 2^n bytes, otherwise narrow bursts are used
	assign M_AXI_ARSIZE	= clogb2((C_M_AXI_DATA_WIDTH/8)-1);
	//INCR burst type is usually used, except for keyhole bursts
	assign M_AXI_ARBURST	= 2'b01;
	assign M_AXI_ARLOCK	= 1'b0;
	//Update value to 4'b0011 if coherent accesses to be used via the Zynq ACP port. Not Allocated, Modifiable, not Bufferable. Not Bufferable since this example is meant to test memory, not intermediate cache.
	assign M_AXI_ARCACHE	= 4'b0010;
	assign M_AXI_ARPROT	= 3'h0;
	assign M_AXI_ARQOS	= 4'h0;
	assign M_AXI_ARVALID	= axi_arvalid;
	//Read and Read Response (R)
	assign M_AXI_RREADY	= axi_rready;
	//Example design I/O
	//Burst size in bytes
	assign burst_size_bytes	= C_M_AXI_BURST_LEN * C_M_AXI_DATA_WIDTH/8;


	//----------------------------
	//Read Address Channel
	//----------------------------

	//The Read Address Channel (AW) provides a similar function to the
	//Write Address channel- to provide the tranfer qualifiers for the burst.

	//In this example, the read address increments in the same
	//manner as the write address channel.

	always @(posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 0) begin
			axi_arvalid <= 1'b0;
		end
		// If previously not valid , start next transaction
		else if (~axi_arvalid && start_single_burst_read) begin
			axi_arvalid <= 1'b1;
		end
		else if (M_AXI_ARREADY && axi_arvalid) begin
			axi_arvalid <= 1'b0;
		end
		else
			axi_arvalid <= axi_arvalid;
	end


	// Next address after ARREADY indicates previous address acceptance
	always @(posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 0) begin
			axi_araddr <= 'b0;
		end
		else if (start_single_burst_read) begin
			if (r_sof)
				axi_araddr <= base_addr;
			else
				axi_araddr <= axi_araddr;
		end
		else if (M_AXI_ARREADY && axi_arvalid) begin
			axi_araddr <= axi_araddr + burst_size_bytes;
		end
		else
			axi_araddr <= axi_araddr;
	end


	//--------------------------------
	//Read Data (and Response) Channel
	//--------------------------------

	 // Forward movement occurs when the channel is valid and ready
	  assign rnext = M_AXI_RVALID && axi_rready;


	// Burst length counter. Uses extra counter register bit to indicate
	// terminal count to reduce decode logic
	always @(posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 0 || start_single_burst_read) begin
			read_index <= 0;
		end
		else if (rnext && (read_index != C_M_AXI_BURST_LEN-1)) begin
			read_index <= read_index + 1;
		end
		else
			read_index <= read_index;
	end


	/*
	 The Read Data channel returns the results of the read request

	 In this example the data checker is always able to accept
	 more data, so no need to throttle the RREADY signal
	 */

	//Flag any read response errors
	assign read_resp_error = axi_rready & M_AXI_RVALID & M_AXI_RRESP[1];


	//--------------------------------
	//Example design throttling
	//--------------------------------

	// For maximum port throughput, this user example code will try to allow
	// each channel to run as independently and as quickly as possible.

	// However, there are times when the flow of data needs to be throtted by
	// the user application. This example application requires that data is
	// not read before it is written and that the write channels do not
	// advance beyond an arbitrary threshold (say to prevent an
	// overrun of the current read address by the write address).

	// From AXI4 Specification, 13.13.1: "If a master requires ordering between
	// read and write transactions, it must ensure that a response is received
	// for the previous transaction before issuing the next transaction."

	// This example accomplishes this user application throttling through:
	// -Reads wait for writes to fully complete
	// -Address writes wait when not read + issued transaction counts pass
	// a parameterized threshold
	// -Writes wait when a not read + active data burst count pass
	// a parameterized threshold

	  //implement master command interface state machine

	always @ ( posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 1'b0 ) begin
			// reset condition
			// All the signals are assigned default values under reset condition
			frame_pulse  <= 1'b0;
		end
		else begin
			// This state is responsible to issue start_single_read pulse to
			// initiate a read transaction. Read transactions will be
			// issued until burst_read_active signal is asserted.
			// read controller
			if (~axi_arvalid && ~burst_read_active && ~frame_pulse) begin
				frame_pulse <= 1'b1;
			end
			else begin
				frame_pulse <= 1'b0; //Negate to generate a pulse
			end
		end
	end //MASTER_EXECUTION_PROC

	always @(posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 1'b0)
			start_single_burst_read <= 1'b0;
		else
			start_single_burst_read <= frame_pulse;
	end

	// burst_read_active signal is asserted when there is a burst write transaction
	// is initiated by the assertion of start_single_burst_write. start_single_burst_read
	// signal remains asserted until the burst read is accepted by the master
	always @(posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 0)
			burst_read_active <= 1'b0;
		//The burst_write_active is asserted when a write burst transaction is initiated
		else if (start_single_burst_read)
			burst_read_active <= 1'b1;
		else if (rnext && M_AXI_RLAST)
			burst_read_active <= 0;
	end

	// Add user logic here

	// User logic ends
	always @(posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 0) begin
			r_img_col_idx <= 0;
			r_img_row_idx <= 0;
		end
		else if (start_single_burst_read
			&& r_img_col_idx == 0
			&& r_img_col_idx == 0) begin
			r_img_col_idx <= C_IMG_WIDTH - C_M_AXI_DATA_WIDTH/8;
			r_img_row_idx <= C_IMG_HEIGHT - 1;
		end
		else if (rnext) begin
			if (r_img_col_idx != 0) begin
				r_img_col_idx <= r_img_col_idx - C_M_AXI_DATA_WIDTH/8;
				r_img_row_idx <= r_img_row_idx;
			end
			else begin
				r_img_col_idx <= C_IMG_WIDTH - C_M_AXI_DATA_WIDTH/8;
				r_img_row_idx <= r_img_row_idx - 1;
			end
		end
		else begin
			r_img_col_idx <= r_img_col_idx;
			r_img_row_idx <= r_img_row_idx;
		end
	end

	always @(posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 0) begin
			r_sof <= 1'b0;
		end
		else if (start_single_burst_read
			&& r_img_col_idx == 0
			&& r_img_col_idx == 0) begin
			r_sof <= 1'b1;
		end
		else if (rnext) begin
			r_sof <= 1'b0;
		end
		else begin
			r_sof <= r_sof;
		end
	end

	always @(posedge M_AXI_ACLK) begin
		if (M_AXI_ARESETN == 0) begin
			r_eol <= 1'b0;
		end
		else if (C_M_AXI_BURST_LEN == 1) begin
			r_eol <= 1'b1;
		end
		else if (rnext) begin
			r_eol <= (r_img_col_idx == C_M_AXI_DATA_WIDTH/8 ? 1'b1 : 1'b0);
		end
		else
			r_eol <= r_eol;
	end

endmodule
